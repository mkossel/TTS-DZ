library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package snn_tts_dataset_pkg is

  -- feature data from the Iris dataset --
  type feature_vector is array (0 to 3) of std_ulogic_vector(0 to 5);
  type feature_array is array (0 to 149) of feature_vector;  
  constant feature_data : feature_array := (
        ( "010111", "001011", "010100", "001010"),  -- (0):   [5.75 2.75 5.   2.5 ]  label: 2   real values: [5.8 2.8 5.1 2.4]
        ( "011000", "001001", "010000", "000100"),  -- (1):   [6.   2.25 4.   1.  ]  label: 1   real values: [6.  2.2 4.  1. ]
        ( "010110", "010001", "000110", "000001"),  -- (2):   [5.5  4.25 1.5  0.25]  label: 0   real values: [5.5 4.2 1.4 0.2]
        ( "011101", "001100", "011001", "000111"),  -- (3):   [7.25 3.   6.25 1.75]  label: 2   real values: [7.3 2.9 6.3 1.8]
        ( "010100", "001110", "000110", "000001"),  -- (4):   [5.   3.5  1.5  0.25]  label: 0   real values: [5.  3.4 1.5 0.2]
        ( "011001", "001101", "011000", "001010"),  -- (5):   [6.25 3.25 6.   2.5 ]  label: 2   real values: [6.3 3.3 6.  2.5]
        ( "010100", "001110", "000101", "000001"),  -- (6):   [5.   3.5  1.25 0.25]  label: 0   real values: [5.  3.5 1.3 0.3]
        ( "011011", "001100", "010011", "000110"),  -- (7):   [6.75 3.   4.75 1.5 ]  label: 1   real values: [6.7 3.1 4.7 1.5]
        ( "011011", "001011", "010011", "000110"),  -- (8):   [6.75 2.75 4.75 1.5 ]  label: 1   real values: [6.8 2.8 4.8 1.4]
        ( "011000", "001011", "010000", "000101"),  -- (9):   [6.   2.75 4.   1.25]  label: 1   real values: [6.1 2.8 4.  1.3]
        ( "011000", "001010", "010110", "000110"),  -- (10):  [6.   2.5  5.5  1.5 ]  label: 2   real values: [6.1 2.6 5.6 1.4]
        ( "011010", "001101", "010010", "000110"),  -- (11):  [6.5  3.25 4.5  1.5 ]  label: 1   real values: [6.4 3.2 4.5 1.5]
        ( "011000", "001011", "010011", "000101"),  -- (12):  [6.   2.75 4.75 1.25]  label: 1   real values: [6.1 2.8 4.7 1.2]
        ( "011010", "001011", "010010", "000110"),  -- (13):  [6.5  2.75 4.5  1.5 ]  label: 1   real values: [6.5 2.8 4.6 1.5]
        ( "011000", "001100", "010011", "000110"),  -- (14):  [6.   3.   4.75 1.5 ]  label: 1   real values: [6.1 2.9 4.7 1.4]
        ( "010100", "001100", "000110", "000000"),  -- (15):  [5.   3.   1.5  0.  ]  label: 0   real values: [4.9 3.1 1.5 0.1]
        ( "011000", "001100", "010010", "000110"),  -- (16):  [6.   3.   4.5  1.5 ]  label: 1   real values: [6.  2.9 4.5 1.5]
        ( "010110", "001010", "010010", "000101"),  -- (17):  [5.5  2.5  4.5  1.25]  label: 1   real values: [5.5 2.6 4.4 1.2]
        ( "010011", "001100", "000110", "000001"),  -- (18):  [4.75 3.   1.5  0.25]  label: 0   real values: [4.8 3.  1.4 0.3]
        ( "010110", "010000", "000101", "000010"),  -- (19):  [5.5  4.   1.25 0.5 ]  label: 0   real values: [5.4 3.9 1.3 0.4]
        ( "010110", "001011", "010100", "001000"),  -- (20):  [5.5  2.75 5.   2.  ]  label: 2   real values: [5.6 2.8 4.9 2. ]
        ( "010110", "001100", "010010", "000110"),  -- (21):  [5.5  3.   4.5  1.5 ]  label: 1   real values: [5.6 3.  4.5 1.5]
        ( "010011", "001110", "001000", "000001"),  -- (22):  [4.75 3.5  2.   0.25]  label: 0   real values: [4.8 3.4 1.9 0.2]
        ( "010010", "001100", "000110", "000001"),  -- (23):  [4.5  3.   1.5  0.25]  label: 0   real values: [4.4 2.9 1.4 0.2]
        ( "011001", "001011", "010011", "000111"),  -- (24):  [6.25 2.75 4.75 1.75]  label: 2   real values: [6.2 2.8 4.8 1.8]
        ( "010010", "001110", "000100", "000001"),  -- (25):  [4.5  3.5  1.   0.25]  label: 0   real values: [4.6 3.6 1.  0.2]
        ( "010100", "001111", "001000", "000010"),  -- (26):  [5.   3.75 2.   0.5 ]  label: 0   real values: [5.1 3.8 1.9 0.4]
        ( "011001", "001100", "010001", "000101"),  -- (27):  [6.25 3.   4.25 1.25]  label: 1   real values: [6.2 2.9 4.3 1.3]
        ( "010100", "001001", "001101", "000100"),  -- (28):  [5.   2.25 3.25 1.  ]  label: 1   real values: [5.  2.3 3.3 1. ]
        ( "010100", "001110", "000110", "000010"),  -- (29):  [5.   3.5  1.5  0.5 ]  label: 0   real values: [5.  3.4 1.6 0.4]
        ( "011010", "001100", "010110", "000111"),  -- (30):  [6.5  3.   5.5  1.75]  label: 2   real values: [6.4 3.1 5.5 1.8]
        ( "010110", "001100", "010010", "000110"),  -- (31):  [5.5  3.   4.5  1.5 ]  label: 1   real values: [5.4 3.  4.5 1.5]
        ( "010101", "001110", "000110", "000001"),  -- (32):  [5.25 3.5  1.5  0.25]  label: 0   real values: [5.2 3.5 1.5 0.2]
        ( "011000", "001100", "010100", "000111"),  -- (33):  [6.   3.   5.   1.75]  label: 2   real values: [6.1 3.  4.9 1.8]
        ( "011010", "001011", "010110", "001001"),  -- (34):  [6.5  2.75 5.5  2.25]  label: 2   real values: [6.4 2.8 5.6 2.2]
        ( "010101", "001011", "010000", "000110"),  -- (35):  [5.25 2.75 4.   1.5 ]  label: 1   real values: [5.2 2.7 3.9 1.4]
        ( "010111", "001111", "000111", "000001"),  -- (36):  [5.75 3.75 1.75 0.25]  label: 0   real values: [5.7 3.8 1.7 0.3]
        ( "011000", "001011", "010100", "000110"),  -- (37):  [6.   2.75 5.   1.5 ]  label: 1   real values: [6.  2.7 5.1 1.6]
        ( "011000", "001100", "010001", "000110"),  -- (38):  [6.   3.   4.25 1.5 ]  label: 1   real values: [5.9 3.  4.2 1.5]
        ( "010111", "001010", "010000", "000101"),  -- (39):  [5.75 2.5  4.   1.25]  label: 1   real values: [5.8 2.6 4.  1.2]
        ( "011011", "001100", "010110", "001000"),  -- (40):  [6.75 3.   5.5  2.  ]  label: 2   real values: [6.8 3.  5.5 2.1]
        ( "010011", "001101", "000101", "000001"),  -- (41):  [4.75 3.25 1.25 0.25]  label: 0   real values: [4.7 3.2 1.3 0.2]
        ( "011100", "001100", "010100", "001001"),  -- (42):  [7.   3.   5.   2.25]  label: 2   real values: [6.9 3.1 5.1 2.3]
        ( "010100", "001110", "000110", "000010"),  -- (43):  [5.   3.5  1.5  0.5 ]  label: 0   real values: [5.  3.5 1.6 0.6]
        ( "010110", "001111", "000110", "000001"),  -- (44):  [5.5  3.75 1.5  0.25]  label: 0   real values: [5.4 3.7 1.5 0.2]
        ( "010100", "001000", "001110", "000100"),  -- (45):  [5.   2.   3.5  1.  ]  label: 1   real values: [5.  2.  3.5 1. ]
        ( "011010", "001100", "010110", "000111"),  -- (46):  [6.5  3.   5.5  1.75]  label: 2   real values: [6.5 3.  5.5 1.8]
        ( "011011", "001101", "010111", "001010"),  -- (47):  [6.75 3.25 5.75 2.5 ]  label: 2   real values: [6.7 3.3 5.7 2.5]
        ( "011000", "001001", "010100", "000110"),  -- (48):  [6.   2.25 5.   1.5 ]  label: 2   real values: [6.  2.2 5.  1.5]
        ( "011011", "001010", "010111", "000111"),  -- (49):  [6.75 2.5  5.75 1.75]  label: 2   real values: [6.7 2.5 5.8 1.8]
        ( "010110", "001010", "010000", "000100"),  -- (50):  [5.5  2.5  4.   1.  ]  label: 1   real values: [5.6 2.5 3.9 1.1]
        ( "011111", "001100", "011000", "001001"),  -- (51):  [7.75 3.   6.   2.25]  label: 2   real values: [7.7 3.  6.1 2.3]
        ( "011001", "001101", "010011", "000110"),  -- (52):  [6.25 3.25 4.75 1.5 ]  label: 1   real values: [6.3 3.3 4.7 1.6]
        ( "010110", "001010", "001111", "000100"),  -- (53):  [5.5  2.5  3.75 1.  ]  label: 1   real values: [5.5 2.4 3.8 1.1]
        ( "011001", "001011", "010100", "000111"),  -- (54):  [6.25 2.75 5.   1.75]  label: 2   real values: [6.3 2.7 4.9 1.8]
        ( "011001", "001011", "010100", "000110"),  -- (55):  [6.25 2.75 5.   1.5 ]  label: 2   real values: [6.3 2.8 5.1 1.5]
        ( "010100", "001010", "010010", "000111"),  -- (56):  [5.   2.5  4.5  1.75]  label: 2   real values: [4.9 2.5 4.5 1.7]
        ( "011001", "001010", "010100", "001000"),  -- (57):  [6.25 2.5  5.   2.  ]  label: 2   real values: [6.3 2.5 5.  1.9]
        ( "011100", "001101", "010011", "000110"),  -- (58):  [7.   3.25 4.75 1.5 ]  label: 1   real values: [7.  3.2 4.7 1.4]
        ( "011010", "001100", "010101", "001000"),  -- (59):  [6.5  3.   5.25 2.  ]  label: 2   real values: [6.5 3.  5.2 2. ]
        ( "011000", "001110", "010010", "000110"),  -- (60):  [6.   3.5  4.5  1.5 ]  label: 1   real values: [6.  3.4 4.5 1.6]
        ( "010011", "001100", "000110", "000001"),  -- (61):  [4.75 3.   1.5  0.25]  label: 0   real values: [4.8 3.1 1.6 0.2]
        ( "010111", "001011", "010100", "001000"),  -- (62):  [5.75 2.75 5.   2.  ]  label: 2   real values: [5.8 2.7 5.1 1.9]
        ( "010110", "001011", "010001", "000101"),  -- (63):  [5.5  2.75 4.25 1.25]  label: 1   real values: [5.6 2.7 4.2 1.3]
        ( "010110", "001100", "001110", "000101"),  -- (64):  [5.5  3.   3.5  1.25]  label: 1   real values: [5.6 2.9 3.6 1.3]
        ( "010110", "001010", "010000", "000101"),  -- (65):  [5.5  2.5  4.   1.25]  label: 1   real values: [5.5 2.5 4.  1.3]
        ( "011000", "001100", "010010", "000110"),  -- (66):  [6.   3.   4.5  1.5 ]  label: 1   real values: [6.1 3.  4.6 1.4]
        ( "011101", "001101", "011000", "000111"),  -- (67):  [7.25 3.25 6.   1.75]  label: 2   real values: [7.2 3.2 6.  1.8]
        ( "010101", "001111", "000110", "000001"),  -- (68):  [5.25 3.75 1.5  0.25]  label: 0   real values: [5.3 3.7 1.5 0.2]
        ( "010001", "001100", "000100", "000000"),  -- (69):  [4.25 3.   1.   0.  ]  label: 0   real values: [4.3 3.  1.1 0.1]
        ( "011010", "001011", "010101", "001000"),  -- (70):  [6.5  2.75 5.25 2.  ]  label: 2   real values: [6.4 2.7 5.3 1.9]
        ( "010111", "001100", "010001", "000101"),  -- (71):  [5.75 3.   4.25 1.25]  label: 1   real values: [5.7 3.  4.2 1.2]
        ( "010110", "001110", "000111", "000001"),  -- (72):  [5.5  3.5  1.75 0.25]  label: 0   real values: [5.4 3.4 1.7 0.2]
        ( "010111", "010010", "000110", "000010"),  -- (73):  [5.75 4.5  1.5  0.5 ]  label: 0   real values: [5.7 4.4 1.5 0.4]
        ( "011100", "001100", "010100", "000110"),  -- (74):  [7.   3.   5.   1.5 ]  label: 1   real values: [6.9 3.1 4.9 1.5]
        ( "010010", "001100", "000110", "000001"),  -- (75):  [4.5  3.   1.5  0.25]  label: 0   real values: [4.6 3.1 1.5 0.2]
        ( "011000", "001100", "010100", "000111"),  -- (76):  [6.   3.   5.   1.75]  label: 2   real values: [5.9 3.  5.1 1.8]
        ( "010100", "001010", "001100", "000100"),  -- (77):  [5.   2.5  3.   1.  ]  label: 1   real values: [5.1 2.5 3.  1.1]
        ( "010010", "001110", "000110", "000001"),  -- (78):  [4.5  3.5  1.5  0.25]  label: 0   real values: [4.6 3.4 1.4 0.3]
        ( "011001", "001001", "010010", "000110"),  -- (79):  [6.25 2.25 4.5  1.5 ]  label: 1   real values: [6.2 2.2 4.5 1.5]
        ( "011101", "001110", "011000", "001010"),  -- (80):  [7.25 3.5  6.   2.5 ]  label: 2   real values: [7.2 3.6 6.1 2.5]
        ( "010111", "001100", "010001", "000101"),  -- (81):  [5.75 3.   4.25 1.25]  label: 1   real values: [5.7 2.9 4.2 1.3]
        ( "010011", "001100", "000110", "000000"),  -- (82):  [4.75 3.   1.5  0.  ]  label: 0   real values: [4.8 3.  1.4 0.1]
        ( "011100", "001100", "011000", "001000"),  -- (83):  [7.   3.   6.   2.  ]  label: 2   real values: [7.1 3.  5.9 2.1]
        ( "011100", "001101", "010111", "001001"),  -- (84):  [7.   3.25 5.75 2.25]  label: 2   real values: [6.9 3.2 5.7 2.3]
        ( "011010", "001100", "010111", "001001"),  -- (85):  [6.5  3.   5.75 2.25]  label: 2   real values: [6.5 3.  5.8 2.2]
        ( "011010", "001011", "010110", "001000"),  -- (86):  [6.5  2.75 5.5  2.  ]  label: 2   real values: [6.4 2.8 5.6 2.1]
        ( "010100", "001111", "000110", "000001"),  -- (87):  [5.   3.75 1.5  0.25]  label: 0   real values: [5.1 3.8 1.6 0.2]
        ( "010011", "001110", "000110", "000001"),  -- (88):  [4.75 3.5  1.5  0.25]  label: 0   real values: [4.8 3.4 1.6 0.2]
        ( "011010", "001101", "010100", "001000"),  -- (89):  [6.5  3.25 5.   2.  ]  label: 2   real values: [6.5 3.2 5.1 2. ]
        ( "011011", "001101", "010111", "001000"),  -- (90):  [6.75 3.25 5.75 2.  ]  label: 2   real values: [6.7 3.3 5.7 2.1]
        ( "010010", "001001", "000101", "000001"),  -- (91):  [4.5  2.25 1.25 0.25]  label: 0   real values: [4.5 2.3 1.3 0.3]
        ( "011001", "001110", "010110", "001001"),  -- (92):  [6.25 3.5  5.5  2.25]  label: 2   real values: [6.2 3.4 5.4 2.3]
        ( "010100", "001100", "000110", "000001"),  -- (93):  [5.   3.   1.5  0.25]  label: 0   real values: [4.9 3.  1.4 0.2]
        ( "010111", "001010", "010100", "001000"),  -- (94):  [5.75 2.5  5.   2.  ]  label: 2   real values: [5.7 2.5 5.  2. ]
        ( "011100", "001100", "010110", "001000"),  -- (95):  [7.   3.   5.5  2.  ]  label: 2   real values: [6.9 3.1 5.4 2.1]
        ( "010010", "001101", "000101", "000001"),  -- (96):  [4.5  3.25 1.25 0.25]  label: 0   real values: [4.4 3.2 1.3 0.2]
        ( "010100", "001110", "000110", "000001"),  -- (97):  [5.   3.5  1.5  0.25]  label: 0   real values: [5.  3.6 1.4 0.2]
        ( "011101", "001100", "010111", "000110"),  -- (98):  [7.25 3.   5.75 1.5 ]  label: 2   real values: [7.2 3.  5.8 1.6]
        ( "010100", "001110", "000110", "000001"),  -- (99):  [5.   3.5  1.5  0.25]  label: 0   real values: [5.1 3.5 1.4 0.3]
        ( "010010", "001100", "000101", "000001"),  -- (100): [4.5  3.   1.25 0.25]  label: 0   real values: [4.4 3.  1.3 0.2]
        ( "010110", "010000", "000111", "000010"),  -- (101): [5.5  4.   1.75 0.5 ]  label: 0   real values: [5.4 3.9 1.7 0.4]
        ( "010110", "001001", "010000", "000101"),  -- (102): [5.5  2.25 4.   1.25]  label: 1   real values: [5.5 2.3 4.  1.3]
        ( "011011", "001101", "011000", "001001"),  -- (103): [6.75 3.25 6.   2.25]  label: 2   real values: [6.8 3.2 5.9 2.3]
        ( "011110", "001100", "011010", "001000"),  -- (104): [7.5  3.   6.5  2.  ]  label: 2   real values: [7.6 3.  6.6 2.1]
        ( "010100", "001110", "000110", "000001"),  -- (105): [5.   3.5  1.5  0.25]  label: 0   real values: [5.1 3.5 1.4 0.2]
        ( "010100", "001100", "000110", "000000"),  -- (106): [5.   3.   1.5  0.  ]  label: 0   real values: [4.9 3.1 1.5 0.1]
        ( "010101", "001110", "000110", "000001"),  -- (107): [5.25 3.5  1.5  0.25]  label: 0   real values: [5.2 3.4 1.4 0.2]
        ( "010111", "001011", "010010", "000101"),  -- (108): [5.75 2.75 4.5  1.25]  label: 1   real values: [5.7 2.8 4.5 1.3]
        ( "011010", "001100", "010010", "000110"),  -- (109): [6.5  3.   4.5  1.5 ]  label: 1   real values: [6.6 3.  4.4 1.4]
        ( "010100", "001101", "000101", "000001"),  -- (110): [5.   3.25 1.25 0.25]  label: 0   real values: [5.  3.2 1.2 0.2]
        ( "010100", "001101", "000111", "000010"),  -- (111): [5.   3.25 1.75 0.5 ]  label: 0   real values: [5.1 3.3 1.7 0.5]
        ( "011010", "001100", "010001", "000101"),  -- (112): [6.5  3.   4.25 1.25]  label: 1   real values: [6.4 2.9 4.3 1.3]
        ( "010110", "001110", "000110", "000010"),  -- (113): [5.5  3.5  1.5  0.5 ]  label: 0   real values: [5.4 3.4 1.5 0.4]
        ( "011111", "001010", "011100", "001001"),  -- (114): [7.75 2.5  7.   2.25]  label: 2   real values: [7.7 2.6 6.9 2.3]
        ( "010100", "001010", "001101", "000100"),  -- (115): [5.   2.5  3.25 1.  ]  label: 1   real values: [4.9 2.4 3.3 1. ]
        ( "011111", "001111", "011010", "001000"),  -- (116): [7.75 3.75 6.5  2.  ]  label: 2   real values: [7.9 3.8 6.4 2. ]
        ( "011011", "001100", "010010", "000110"),  -- (117): [6.75 3.   4.5  1.5 ]  label: 1   real values: [6.7 3.1 4.4 1.4]
        ( "010101", "010000", "000110", "000000"),  -- (118): [5.25 4.   1.5  0.  ]  label: 0   real values: [5.2 4.1 1.5 0.1]
        ( "011000", "001100", "010011", "000111"),  -- (119): [6.   3.   4.75 1.75]  label: 2   real values: [6.  3.  4.8 1.8]
        ( "010111", "010000", "000101", "000001"),  -- (120): [5.75 4.   1.25 0.25]  label: 0   real values: [5.8 4.  1.2 0.2]
        ( "011111", "001011", "011011", "001000"),  -- (121): [7.75 2.75 6.75 2.  ]  label: 2   real values: [7.7 2.8 6.7 2. ]
        ( "010100", "001111", "000110", "000001"),  -- (122): [5.   3.75 1.5  0.25]  label: 0   real values: [5.1 3.8 1.5 0.3]
        ( "010011", "001101", "000110", "000001"),  -- (123): [4.75 3.25 1.5  0.25]  label: 0   real values: [4.7 3.2 1.6 0.2]
        ( "011110", "001011", "011000", "001000"),  -- (124): [7.5  2.75 6.   2.  ]  label: 2   real values: [7.4 2.8 6.1 1.9]
        ( "010100", "001101", "000110", "000001"),  -- (125): [5.   3.25 1.5  0.25]  label: 0   real values: [5.  3.3 1.4 0.2]
        ( "011001", "001110", "010110", "001010"),  -- (126): [6.25 3.5  5.5  2.5 ]  label: 2   real values: [6.3 3.4 5.6 2.4]
        ( "010111", "001011", "010000", "000101"),  -- (127): [5.75 2.75 4.   1.25]  label: 1   real values: [5.7 2.8 4.1 1.3]
        ( "010111", "001011", "010000", "000101"),  -- (128): [5.75 2.75 4.   1.25]  label: 1   real values: [5.8 2.7 3.9 1.2]
        ( "010111", "001010", "001110", "000100"),  -- (129): [5.75 2.5  3.5  1.  ]  label: 1   real values: [5.7 2.6 3.5 1. ]
        ( "011010", "001101", "010101", "001001"),  -- (130): [6.5  3.25 5.25 2.25]  label: 2   real values: [6.4 3.2 5.3 2.3]
        ( "011011", "001100", "010101", "001001"),  -- (131): [6.75 3.   5.25 2.25]  label: 2   real values: [6.7 3.  5.2 2.3]
        ( "011001", "001010", "010100", "000110"),  -- (132): [6.25 2.5  5.   1.5 ]  label: 1   real values: [6.3 2.5 4.9 1.5]
        ( "011011", "001100", "010100", "000111"),  -- (133): [6.75 3.   5.   1.75]  label: 1   real values: [6.7 3.  5.  1.7]
        ( "010100", "001100", "000110", "000001"),  -- (134): [5.   3.   1.5  0.25]  label: 0   real values: [5.  3.  1.6 0.2]
        ( "010110", "001010", "001111", "000100"),  -- (135): [5.5  2.5  3.75 1.  ]  label: 1   real values: [5.5 2.4 3.7 1. ]
        ( "011011", "001100", "010110", "001010"),  -- (136): [6.75 3.   5.5  2.5 ]  label: 2   real values: [6.7 3.1 5.6 2.4]
        ( "010111", "001011", "010100", "001000"),  -- (137): [5.75 2.75 5.   2.  ]  label: 2   real values: [5.8 2.7 5.1 1.9]
        ( "010100", "001110", "000110", "000001"),  -- (138): [5.   3.5  1.5  0.25]  label: 0   real values: [5.1 3.4 1.5 0.2]
        ( "011010", "001100", "010010", "000101"),  -- (139): [6.5  3.   4.5  1.25]  label: 1   real values: [6.6 2.9 4.6 1.3]
        ( "010110", "001100", "010000", "000101"),  -- (140): [5.5  3.   4.   1.25]  label: 1   real values: [5.6 3.  4.1 1.3]
        ( "011000", "001101", "010011", "000111"),  -- (141): [6.   3.25 4.75 1.75]  label: 1   real values: [5.9 3.2 4.8 1.8]
        ( "011001", "001001", "010010", "000101"),  -- (142): [6.25 2.25 4.5  1.25]  label: 1   real values: [6.3 2.3 4.4 1.3]
        ( "010110", "001110", "000101", "000001"),  -- (143): [5.5  3.5  1.25 0.25]  label: 0   real values: [5.5 3.5 1.3 0.2]
        ( "010100", "001111", "000110", "000010"),  -- (144): [5.   3.75 1.5  0.5 ]  label: 0   real values: [5.1 3.7 1.5 0.4]
        ( "010100", "001100", "000110", "000000"),  -- (145): [5.   3.   1.5  0.  ]  label: 0   real values: [4.9 3.1 1.5 0.1]
        ( "011001", "001100", "010110", "000111"),  -- (146): [6.25 3.   5.5  1.75]  label: 2   real values: [6.3 2.9 5.6 1.8]
        ( "010111", "001011", "010000", "000100"),  -- (147): [5.75 2.75 4.   1.  ]  label: 1   real values: [5.8 2.7 4.1 1. ]
        ( "011111", "001111", "011011", "001001"),  -- (148): [7.75 3.75 6.75 2.25]  label: 2   real values: [7.7 3.8 6.7 2.2]
        ( "010010", "001101", "000110", "000001")   -- (149): [4.5  3.25 1.5  0.25]  label: 0   real values: [4.6 3.2 1.4 0.2]		
        );
	
  type feature_label is array (0 to 149) of integer;  
  constant feature_label_value : feature_label := (
	2,
	1,
	0,
	2,
	0,
	2,
	0,
	1,
	1,
	1,
	2,
	1,
	1,
	1,
	1,
	0,
	1,
	1,
	0,
	0,
	2,
	1,
	0,
	0,
	2,
	0,
	0,
	1,
	1,
	0,
	2,
	1,
	0,
	2,
	2,
	1,
	0,
	1,
	1,
	1,
	2,
	0,
	2,
	0,
	0,
	1,
	2,
	2,
	2,
	2,
	1,
	2,
	1,
	1,
	2,
	2,
	2,
	2,
	1,
	2,
	1,
	0,
	2,
	1,
	1,
	1,
	1,
	2,
	0,
	0,
	2,
	1,
	0,
	0,
	1,
	0,
	2,
	1,
	0,
	1,
	2,
	1,
	0,
	2,
	2,
	2,
	2,
	0,
	0,
	2,
	2,
	0,
	2,
	0,
	2,
	2,
	0,
	0,
	2,
	0,
	0,
	0,
	1,
	2,
	2,
	0,
	0,
	0,
	1,
	1,
	0,
	0,
	1,
	0,
	2,
	1,
	2,
	1,
	0,
	2,
	0,
	2,
	0,
	0,
	2,
	0,
	2,
	1,
	1,
	1,
	2,
	2,
	1,
	1,
	0,
	1,
	2,
	2,
	0,
	1,
	1,
	1,
	1,
	0,
	0,
	0,
	2,
	1,
	2,
	0	
	);
  
end package snn_tts_dataset_pkg;


package body snn_tts_dataset_pkg is



end package body snn_tts_dataset_pkg;
